VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO top_tukka_proj
  CLASS BLOCK ;
  FOREIGN top_tukka_proj ;
  ORIGIN 0.000 0.000 ;
  SIZE 1500.000 BY 1500.000 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT -0.880 8.080 0.720 1489.360 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -0.880 8.080 1500.560 9.680 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -0.880 1487.760 1500.560 1489.360 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1498.960 8.080 1500.560 1489.360 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 22.240 4.780 23.840 1492.660 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 175.840 4.780 177.440 1492.660 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 329.440 4.780 331.040 1492.660 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 483.040 4.780 484.640 1492.660 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 636.640 4.780 638.240 1492.660 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 790.240 4.780 791.840 1492.660 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 943.840 4.780 945.440 1492.660 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1097.440 4.780 1099.040 1492.660 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1251.040 4.780 1252.640 1492.660 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1404.640 4.780 1406.240 1492.660 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -4.180 31.530 1503.860 33.130 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -4.180 184.710 1503.860 186.310 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -4.180 337.890 1503.860 339.490 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -4.180 491.070 1503.860 492.670 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -4.180 644.250 1503.860 645.850 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -4.180 797.430 1503.860 799.030 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -4.180 950.610 1503.860 952.210 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -4.180 1103.790 1503.860 1105.390 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -4.180 1256.970 1503.860 1258.570 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -4.180 1410.150 1503.860 1411.750 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT -4.180 4.780 -2.580 1492.660 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -4.180 4.780 1503.860 6.380 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -4.180 1491.060 1503.860 1492.660 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1502.260 4.780 1503.860 1492.660 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 25.540 4.780 27.140 1492.660 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 179.140 4.780 180.740 1492.660 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 332.740 4.780 334.340 1492.660 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 486.340 4.780 487.940 1492.660 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 639.940 4.780 641.540 1492.660 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 793.540 4.780 795.140 1492.660 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 947.140 4.780 948.740 1492.660 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1100.740 4.780 1102.340 1492.660 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1254.340 4.780 1255.940 1492.660 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1407.940 4.780 1409.540 1492.660 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -4.180 34.830 1503.860 36.430 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -4.180 188.010 1503.860 189.610 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -4.180 341.190 1503.860 342.790 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -4.180 494.370 1503.860 495.970 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -4.180 647.550 1503.860 649.150 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -4.180 800.730 1503.860 802.330 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -4.180 953.910 1503.860 955.510 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -4.180 1107.090 1503.860 1108.690 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -4.180 1260.270 1503.860 1261.870 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -4.180 1413.450 1503.860 1415.050 ;
    END
  END VSS
  PIN address[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1496.000 1159.200 1499.000 1159.760 ;
    END
  END address[0]
  PIN address[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 853.440 1496.000 854.000 1499.000 ;
    END
  END address[1]
  PIN address[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 910.560 4.000 911.120 ;
    END
  END address[2]
  PIN address[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 302.400 1.000 302.960 4.000 ;
    END
  END address[3]
  PIN address[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1496.000 396.480 1499.000 397.040 ;
    END
  END address[4]
  PIN address[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 379.680 4.000 380.240 ;
    END
  END address[5]
  PIN address[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1216.320 1.000 1216.880 4.000 ;
    END
  END address[6]
  PIN address[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 225.120 4.000 225.680 ;
    END
  END address[7]
  PIN clk1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 151.200 4.000 151.760 ;
    END
  END clk1
  PIN clk2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1496.000 473.760 1499.000 474.320 ;
    END
  END clk2
  PIN cs
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 1216.320 4.000 1216.880 ;
    END
  END cs
  PIN error
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 608.160 4.000 608.720 ;
    END
  END error
  PIN read_data[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1444.800 1.000 1445.360 4.000 ;
    END
  END read_data[0]
  PIN read_data[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 1061.760 4.000 1062.320 ;
    END
  END read_data[10]
  PIN read_data[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 16.800 1496.000 17.360 1499.000 ;
    END
  END read_data[11]
  PIN read_data[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 759.360 4.000 759.920 ;
    END
  END read_data[12]
  PIN read_data[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 930.720 1496.000 931.280 1499.000 ;
    END
  END read_data[13]
  PIN read_data[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1496.000 322.560 1499.000 323.120 ;
    END
  END read_data[14]
  PIN read_data[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 1139.040 4.000 1139.600 ;
    END
  END read_data[15]
  PIN read_data[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1496.000 551.040 1499.000 551.600 ;
    END
  END read_data[16]
  PIN read_data[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1387.680 1496.000 1388.240 1499.000 ;
    END
  END read_data[17]
  PIN read_data[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1496.000 1081.920 1499.000 1082.480 ;
    END
  END read_data[18]
  PIN read_data[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 302.400 4.000 302.960 ;
    END
  END read_data[19]
  PIN read_data[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1496.000 1387.680 1499.000 1388.240 ;
    END
  END read_data[1]
  PIN read_data[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1496.000 930.720 1499.000 931.280 ;
    END
  END read_data[20]
  PIN read_data[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 473.760 1496.000 474.320 1499.000 ;
    END
  END read_data[21]
  PIN read_data[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1496.000 1233.120 1499.000 1233.680 ;
    END
  END read_data[22]
  PIN read_data[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1290.240 1.000 1290.800 4.000 ;
    END
  END read_data[23]
  PIN read_data[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1496.000 168.000 1499.000 168.560 ;
    END
  END read_data[24]
  PIN read_data[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 151.200 1.000 151.760 4.000 ;
    END
  END read_data[25]
  PIN read_data[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1004.640 1496.000 1005.200 1499.000 ;
    END
  END read_data[26]
  PIN read_data[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 530.880 1.000 531.440 4.000 ;
    END
  END read_data[27]
  PIN read_data[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 910.560 1.000 911.120 4.000 ;
    END
  END read_data[28]
  PIN read_data[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1496.000 1004.640 1499.000 1005.200 ;
    END
  END read_data[29]
  PIN read_data[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 833.280 4.000 833.840 ;
    END
  END read_data[2]
  PIN read_data[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 94.080 1496.000 94.640 1499.000 ;
    END
  END read_data[30]
  PIN read_data[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 379.680 1.000 380.240 4.000 ;
    END
  END read_data[31]
  PIN read_data[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1139.040 1.000 1139.600 4.000 ;
    END
  END read_data[3]
  PIN read_data[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1159.200 1496.000 1159.760 1499.000 ;
    END
  END read_data[4]
  PIN read_data[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1496.000 16.800 1499.000 17.360 ;
    END
  END read_data[5]
  PIN read_data[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 551.040 1496.000 551.600 1499.000 ;
    END
  END read_data[6]
  PIN read_data[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 1444.800 4.000 1445.360 ;
    END
  END read_data[7]
  PIN read_data[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1367.520 1.000 1368.080 4.000 ;
    END
  END read_data[8]
  PIN read_data[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 624.960 1496.000 625.520 1499.000 ;
    END
  END read_data[9]
  PIN reset_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1496.000 245.280 1499.000 245.840 ;
    END
  END reset_n
  PIN sel_clk2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1496.000 624.960 1499.000 625.520 ;
    END
  END sel_clk2
  PIN we
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1061.760 1.000 1062.320 4.000 ;
    END
  END we
  PIN write_data[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 73.920 4.000 74.480 ;
    END
  END write_data[0]
  PIN write_data[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 1367.520 4.000 1368.080 ;
    END
  END write_data[10]
  PIN write_data[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 776.160 1496.000 776.720 1499.000 ;
    END
  END write_data[11]
  PIN write_data[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 682.080 1.000 682.640 4.000 ;
    END
  END write_data[12]
  PIN write_data[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1.000 0.560 4.000 ;
    END
  END write_data[13]
  PIN write_data[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 682.080 4.000 682.640 ;
    END
  END write_data[14]
  PIN write_data[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 702.240 1496.000 702.800 1499.000 ;
    END
  END write_data[15]
  PIN write_data[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1081.920 1496.000 1082.480 1499.000 ;
    END
  END write_data[16]
  PIN write_data[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1461.600 1496.000 1462.160 1499.000 ;
    END
  END write_data[17]
  PIN write_data[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 322.560 1496.000 323.120 1499.000 ;
    END
  END write_data[18]
  PIN write_data[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 987.840 4.000 988.400 ;
    END
  END write_data[19]
  PIN write_data[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 73.920 1.000 74.480 4.000 ;
    END
  END write_data[1]
  PIN write_data[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1496.000 1461.600 1499.000 1462.160 ;
    END
  END write_data[20]
  PIN write_data[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 530.880 4.000 531.440 ;
    END
  END write_data[21]
  PIN write_data[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 608.160 1.000 608.720 4.000 ;
    END
  END write_data[22]
  PIN write_data[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1496.000 1310.400 1499.000 1310.960 ;
    END
  END write_data[23]
  PIN write_data[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1496.000 94.080 1499.000 94.640 ;
    END
  END write_data[24]
  PIN write_data[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 245.280 1496.000 245.840 1499.000 ;
    END
  END write_data[25]
  PIN write_data[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1496.000 776.160 1499.000 776.720 ;
    END
  END write_data[26]
  PIN write_data[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 225.120 1.000 225.680 4.000 ;
    END
  END write_data[27]
  PIN write_data[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 453.600 1.000 454.160 4.000 ;
    END
  END write_data[28]
  PIN write_data[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 759.360 1.000 759.920 4.000 ;
    END
  END write_data[29]
  PIN write_data[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1496.000 853.440 1499.000 854.000 ;
    END
  END write_data[2]
  PIN write_data[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 833.280 1.000 833.840 4.000 ;
    END
  END write_data[30]
  PIN write_data[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1310.400 1496.000 1310.960 1499.000 ;
    END
  END write_data[31]
  PIN write_data[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1233.120 1496.000 1233.680 1499.000 ;
    END
  END write_data[3]
  PIN write_data[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 168.000 1496.000 168.560 1499.000 ;
    END
  END write_data[4]
  PIN write_data[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 396.480 1496.000 397.040 1499.000 ;
    END
  END write_data[5]
  PIN write_data[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 987.840 1.000 988.400 4.000 ;
    END
  END write_data[6]
  PIN write_data[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 453.600 4.000 454.160 ;
    END
  END write_data[7]
  PIN write_data[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 1290.240 4.000 1290.800 ;
    END
  END write_data[8]
  PIN write_data[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1496.000 702.240 1499.000 702.800 ;
    END
  END write_data[9]
  OBS
      LAYER Metal1 ;
        RECT 6.720 15.380 1492.960 1482.730 ;
      LAYER Metal2 ;
        RECT 0.140 1495.700 16.500 1496.000 ;
        RECT 17.660 1495.700 93.780 1496.000 ;
        RECT 94.940 1495.700 167.700 1496.000 ;
        RECT 168.860 1495.700 244.980 1496.000 ;
        RECT 246.140 1495.700 322.260 1496.000 ;
        RECT 323.420 1495.700 396.180 1496.000 ;
        RECT 397.340 1495.700 473.460 1496.000 ;
        RECT 474.620 1495.700 550.740 1496.000 ;
        RECT 551.900 1495.700 624.660 1496.000 ;
        RECT 625.820 1495.700 701.940 1496.000 ;
        RECT 703.100 1495.700 775.860 1496.000 ;
        RECT 777.020 1495.700 853.140 1496.000 ;
        RECT 854.300 1495.700 930.420 1496.000 ;
        RECT 931.580 1495.700 1004.340 1496.000 ;
        RECT 1005.500 1495.700 1081.620 1496.000 ;
        RECT 1082.780 1495.700 1158.900 1496.000 ;
        RECT 1160.060 1495.700 1232.820 1496.000 ;
        RECT 1233.980 1495.700 1310.100 1496.000 ;
        RECT 1311.260 1495.700 1387.380 1496.000 ;
        RECT 1388.540 1495.700 1461.300 1496.000 ;
        RECT 1462.460 1495.700 1491.140 1496.000 ;
        RECT 0.140 4.300 1491.140 1495.700 ;
        RECT 0.860 4.000 73.620 4.300 ;
        RECT 74.780 4.000 150.900 4.300 ;
        RECT 152.060 4.000 224.820 4.300 ;
        RECT 225.980 4.000 302.100 4.300 ;
        RECT 303.260 4.000 379.380 4.300 ;
        RECT 380.540 4.000 453.300 4.300 ;
        RECT 454.460 4.000 530.580 4.300 ;
        RECT 531.740 4.000 607.860 4.300 ;
        RECT 609.020 4.000 681.780 4.300 ;
        RECT 682.940 4.000 759.060 4.300 ;
        RECT 760.220 4.000 832.980 4.300 ;
        RECT 834.140 4.000 910.260 4.300 ;
        RECT 911.420 4.000 987.540 4.300 ;
        RECT 988.700 4.000 1061.460 4.300 ;
        RECT 1062.620 4.000 1138.740 4.300 ;
        RECT 1139.900 4.000 1216.020 4.300 ;
        RECT 1217.180 4.000 1289.940 4.300 ;
        RECT 1291.100 4.000 1367.220 4.300 ;
        RECT 1368.380 4.000 1444.500 4.300 ;
        RECT 1445.660 4.000 1491.140 4.300 ;
      LAYER Metal3 ;
        RECT 0.090 1462.460 1496.000 1481.900 ;
        RECT 0.090 1461.300 1495.700 1462.460 ;
        RECT 0.090 1445.660 1496.000 1461.300 ;
        RECT 0.090 1444.500 0.700 1445.660 ;
        RECT 4.300 1444.500 1496.000 1445.660 ;
        RECT 0.090 1388.540 1496.000 1444.500 ;
        RECT 0.090 1387.380 1495.700 1388.540 ;
        RECT 0.090 1368.380 1496.000 1387.380 ;
        RECT 0.090 1367.220 0.700 1368.380 ;
        RECT 4.300 1367.220 1496.000 1368.380 ;
        RECT 0.090 1311.260 1496.000 1367.220 ;
        RECT 0.090 1310.100 1495.700 1311.260 ;
        RECT 0.090 1291.100 1496.000 1310.100 ;
        RECT 0.090 1289.940 0.700 1291.100 ;
        RECT 4.300 1289.940 1496.000 1291.100 ;
        RECT 0.090 1233.980 1496.000 1289.940 ;
        RECT 0.090 1232.820 1495.700 1233.980 ;
        RECT 0.090 1217.180 1496.000 1232.820 ;
        RECT 0.090 1216.020 0.700 1217.180 ;
        RECT 4.300 1216.020 1496.000 1217.180 ;
        RECT 0.090 1160.060 1496.000 1216.020 ;
        RECT 0.090 1158.900 1495.700 1160.060 ;
        RECT 0.090 1139.900 1496.000 1158.900 ;
        RECT 0.090 1138.740 0.700 1139.900 ;
        RECT 4.300 1138.740 1496.000 1139.900 ;
        RECT 0.090 1082.780 1496.000 1138.740 ;
        RECT 0.090 1081.620 1495.700 1082.780 ;
        RECT 0.090 1062.620 1496.000 1081.620 ;
        RECT 0.090 1061.460 0.700 1062.620 ;
        RECT 4.300 1061.460 1496.000 1062.620 ;
        RECT 0.090 1005.500 1496.000 1061.460 ;
        RECT 0.090 1004.340 1495.700 1005.500 ;
        RECT 0.090 988.700 1496.000 1004.340 ;
        RECT 0.090 987.540 0.700 988.700 ;
        RECT 4.300 987.540 1496.000 988.700 ;
        RECT 0.090 931.580 1496.000 987.540 ;
        RECT 0.090 930.420 1495.700 931.580 ;
        RECT 0.090 911.420 1496.000 930.420 ;
        RECT 0.090 910.260 0.700 911.420 ;
        RECT 4.300 910.260 1496.000 911.420 ;
        RECT 0.090 854.300 1496.000 910.260 ;
        RECT 0.090 853.140 1495.700 854.300 ;
        RECT 0.090 834.140 1496.000 853.140 ;
        RECT 0.090 832.980 0.700 834.140 ;
        RECT 4.300 832.980 1496.000 834.140 ;
        RECT 0.090 777.020 1496.000 832.980 ;
        RECT 0.090 775.860 1495.700 777.020 ;
        RECT 0.090 760.220 1496.000 775.860 ;
        RECT 0.090 759.060 0.700 760.220 ;
        RECT 4.300 759.060 1496.000 760.220 ;
        RECT 0.090 703.100 1496.000 759.060 ;
        RECT 0.090 701.940 1495.700 703.100 ;
        RECT 0.090 682.940 1496.000 701.940 ;
        RECT 0.090 681.780 0.700 682.940 ;
        RECT 4.300 681.780 1496.000 682.940 ;
        RECT 0.090 625.820 1496.000 681.780 ;
        RECT 0.090 624.660 1495.700 625.820 ;
        RECT 0.090 609.020 1496.000 624.660 ;
        RECT 0.090 607.860 0.700 609.020 ;
        RECT 4.300 607.860 1496.000 609.020 ;
        RECT 0.090 551.900 1496.000 607.860 ;
        RECT 0.090 550.740 1495.700 551.900 ;
        RECT 0.090 531.740 1496.000 550.740 ;
        RECT 0.090 530.580 0.700 531.740 ;
        RECT 4.300 530.580 1496.000 531.740 ;
        RECT 0.090 474.620 1496.000 530.580 ;
        RECT 0.090 473.460 1495.700 474.620 ;
        RECT 0.090 454.460 1496.000 473.460 ;
        RECT 0.090 453.300 0.700 454.460 ;
        RECT 4.300 453.300 1496.000 454.460 ;
        RECT 0.090 397.340 1496.000 453.300 ;
        RECT 0.090 396.180 1495.700 397.340 ;
        RECT 0.090 380.540 1496.000 396.180 ;
        RECT 0.090 379.380 0.700 380.540 ;
        RECT 4.300 379.380 1496.000 380.540 ;
        RECT 0.090 323.420 1496.000 379.380 ;
        RECT 0.090 322.260 1495.700 323.420 ;
        RECT 0.090 303.260 1496.000 322.260 ;
        RECT 0.090 302.100 0.700 303.260 ;
        RECT 4.300 302.100 1496.000 303.260 ;
        RECT 0.090 246.140 1496.000 302.100 ;
        RECT 0.090 244.980 1495.700 246.140 ;
        RECT 0.090 225.980 1496.000 244.980 ;
        RECT 0.090 224.820 0.700 225.980 ;
        RECT 4.300 224.820 1496.000 225.980 ;
        RECT 0.090 168.860 1496.000 224.820 ;
        RECT 0.090 167.700 1495.700 168.860 ;
        RECT 0.090 152.060 1496.000 167.700 ;
        RECT 0.090 150.900 0.700 152.060 ;
        RECT 4.300 150.900 1496.000 152.060 ;
        RECT 0.090 94.940 1496.000 150.900 ;
        RECT 0.090 93.780 1495.700 94.940 ;
        RECT 0.090 74.780 1496.000 93.780 ;
        RECT 0.090 73.620 0.700 74.780 ;
        RECT 4.300 73.620 1496.000 74.780 ;
        RECT 0.090 17.660 1496.000 73.620 ;
        RECT 0.090 16.500 1495.700 17.660 ;
        RECT 0.090 14.700 1496.000 16.500 ;
      LAYER Metal4 ;
        RECT 18.060 14.650 21.940 1481.110 ;
        RECT 24.140 14.650 25.240 1481.110 ;
        RECT 27.440 14.650 175.540 1481.110 ;
        RECT 177.740 14.650 178.840 1481.110 ;
        RECT 181.040 14.650 329.140 1481.110 ;
        RECT 331.340 14.650 332.440 1481.110 ;
        RECT 334.640 14.650 482.740 1481.110 ;
        RECT 484.940 14.650 486.040 1481.110 ;
        RECT 488.240 14.650 636.340 1481.110 ;
        RECT 638.540 14.650 639.640 1481.110 ;
        RECT 641.840 14.650 789.940 1481.110 ;
        RECT 792.140 14.650 793.240 1481.110 ;
        RECT 795.440 14.650 943.540 1481.110 ;
        RECT 945.740 14.650 946.840 1481.110 ;
        RECT 949.040 14.650 1097.140 1481.110 ;
        RECT 1099.340 14.650 1100.440 1481.110 ;
        RECT 1102.640 14.650 1250.740 1481.110 ;
        RECT 1252.940 14.650 1254.040 1481.110 ;
        RECT 1256.240 14.650 1404.340 1481.110 ;
        RECT 1406.540 14.650 1407.640 1481.110 ;
        RECT 1409.840 14.650 1475.460 1481.110 ;
      LAYER Metal5 ;
        RECT 17.980 1109.190 1474.980 1186.020 ;
        RECT 17.980 1105.890 1474.980 1106.590 ;
        RECT 17.980 956.010 1474.980 1103.290 ;
        RECT 17.980 952.710 1474.980 953.410 ;
        RECT 17.980 802.830 1474.980 950.110 ;
        RECT 17.980 799.530 1474.980 800.230 ;
        RECT 17.980 649.650 1474.980 796.930 ;
        RECT 17.980 646.350 1474.980 647.050 ;
        RECT 17.980 496.470 1474.980 643.750 ;
        RECT 17.980 493.170 1474.980 493.870 ;
        RECT 17.980 394.300 1474.980 490.570 ;
  END
END top_tukka_proj
END LIBRARY

